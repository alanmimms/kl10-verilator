`timescale 1ns/1ps
// M8534 CCW
module ccw();
endmodule // ccw

