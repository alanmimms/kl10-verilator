`timescale 1ns/1ps
module cha();
endmodule // cha
