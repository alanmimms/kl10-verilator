`timescale 1ns/1ps
// M8521 CHD
module chd();
endmodule // chd
